// 4-Bit Ripple Carry Adder
// Written by Cole Garrett Shoemaker




module four_bit_RCA (A, B, Cin, S, Cout);
  input [3:0] A, B;
  input Cin;
  output [3:0] S;
  output Cout;

  
  
